LIBRARY IEEE;
LIBRARY ALTERA_MF;
LIBRARY LPM;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ALTERA_MF.ALTERA_MF_COMPONENTS.ALL;
USE LPM.LPM_COMPONENTS.ALL;


ENTITY SRAM IS
	PORT(
		CLOCK          : IN    STD_LOGIC;
		RESETN         : IN    STD_LOGIC;
		IO_WRITE       : IN    STD_LOGIC;
		SRAM_ADHI_EN   : IN    STD_LOGIC;
		SRAM_ADLOW_EN  : IN    STD_LOGIC;
		SRAM_DATA_EN   : IN    STD_LOGIC;
		IO_DATA        : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		SRAM_ADDR      : OUT   STD_LOGIC_VECTOR(17 DOWNTO 0);
		SRAM_OE_N      : OUT   STD_LOGIC;
		SRAM_DQ        : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		SRAM_WE_N      : OUT   STD_LOGIC;
		SRAM_UB_N      : OUT   STD_LOGIC;
		SRAM_LB_N      : OUT   STD_LOGIC;
		SRAM_CE_N      : OUT   STD_LOGIC
	);
END SRAM;

ARCHITECTURE a of SRAM IS
  TYPE STATE_TYPE IS (
	IDLE, SET_HIGH, SET_LOW, GET_DATA, READ_DATA, WRITE1, WRITE2
  );
  SIGNAL STATE     : STATE_TYPE;
  SIGNAL SRAM_DATA : STD_LOGIC_VECTOR(15 DOWNTO 0);
  SIGNAL SRAM_MODE : STD_LOGIC_VECTOR(3 DOWNTO 0);
  BEGIN
    PROCESS(CLOCK, RESETN)
      BEGIN
        IF RESETN = '0' THEN
          STATE <= IDLE;
        ELSIF (RISING_EDGE(CLOCK)) THEN
		  CASE STATE IS
            WHEN IDLE =>
              SRAM_WE_N <= '1';
              IO_DATA   <= "ZZZZZZZZZZZZZZZZ";
			  CASE SRAM_MODE IS
				WHEN "1100" => STATE <= SET_HIGH;
				WHEN "1010" => STATE <= SET_LOW;
				WHEN "0001" => STATE <= READ_DATA;
				WHEN "1001" => STATE <= WRITE1;
				WHEN OTHERS => STATE <= IDLE;
			  END CASE;
			WHEN SET_HIGH =>
			  SRAM_ADDR(17 DOWNTO 16) <= IO_DATA(1 DOWNTO 0);
			  CASE SRAM_MODE IS
				WHEN "1100" => STATE <= SET_HIGH;
				WHEN OTHERS => STATE <= GET_DATA;
			  END CASE;
			WHEN SET_LOW =>
			  SRAM_ADDR(15 DOWNTO 0) <= IO_DATA(15 DOWNTO 0);
			  CASE SRAM_MODE IS
				WHEN "1010" => STATE <= SET_HIGH;
				WHEN OTHERS => STATE <= GET_DATA;
			  END CASE;
			WHEN GET_DATA =>
			  SRAM_DATA <= SRAM_DQ;
			  STATE <= IDLE;
			WHEN READ_DATA =>
			  IO_DATA <= SRAM_DATA;
			  CASE SRAM_MODE IS
				WHEN "0001" => STATE <= READ_DATA;
				WHEN OTHERS => STATE <= IDLE;
			  END CASE;
			WHEN WRITE1 =>
			  SRAM_DATA <= IO_DATA;
			  SRAM_DQ   <= SRAM_DATA;
			  CASE SRAM_MODE IS
				WHEN "1001" => STATE <= WRITE1;
				WHEN OTHERS => STATE <= WRITE2;
			  END CASE;
			WHEN WRITE2 =>
			  SRAM_WE_N <= '0';
			  SRAM_DQ   <= SRAM_DATA;
			  STATE <= IDLE;
			WHEN OTHERS =>
			  STATE <=IDLE;
          END CASE;
        END IF;
      END PROCESS;
    --Combined Mode Vector  
    SRAM_MODE <= IO_WRITE & SRAM_ADHI_EN & SRAM_ADLOW_EN & SRAM_DATA_EN;
    --Constants
    SRAM_CE_N <= '0';
    SRAM_UB_N <= '0';
	SRAM_LB_N <= '0';
	--Always avaliable read unless WE is active
	SRAM_OE_N <= '0';
	

  END a;
