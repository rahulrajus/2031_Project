LIBRARY IEEE;
LIBRARY ALTERA_MF;
LIBRARY LPM;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE ALTERA_MF.ALTERA_MF_COMPONENTS.ALL;
USE LPM.LPM_COMPONENTS.ALL;


ENTITY SRAM IS
	PORT(
		CLOCK          : IN    STD_LOGIC;
		RESETN         : IN    STD_LOGIC;
		IO_WRITE       : IN    STD_LOGIC;
		SRAM_ADHI_EN   : IN    STD_LOGIC;
		SRAM_ADLOW_EN  : IN    STD_LOGIC;
		SRAM_DATA_EN   : IN    STD_LOGIC;
		IO_CYCLE       : IN    STD_LOGIC;
		IO_DATA        : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		SRAM_ADDR      : OUT   STD_LOGIC_VECTOR(17 DOWNTO 0);
		SRAM_OE_N      : OUT   STD_LOGIC;
		SRAM_DQ        : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		SRAM_WE_N      : OUT   STD_LOGIC;
		SRAM_UB_N      : OUT   STD_LOGIC;
		SRAM_LB_N      : OUT   STD_LOGIC;
		SRAM_CE_N      : OUT   STD_LOGIC
	);
END SRAM;

ARCHITECTURE a of SRAM IS
  TYPE STATE_TYPE IS (
	IDLE, WRITE_DATA, WRITE_DATA2, SET_HIGH, SET_LOW
  );
  SIGNAL STATE       : STATE_TYPE;
  SIGNAL SRAM_DATA   : STD_LOGIC_VECTOR(15 DOWNTO 0);
  SIGNAL SRAM_MODE   : STD_LOGIC_VECTOR(3 DOWNTO 0);
  SIGNAL IO_DATA_INT : STD_LOGIC;
  
  BEGIN
	--Combined Mode Vector  
    SRAM_MODE <= IO_WRITE & SRAM_ADHI_EN & SRAM_ADLOW_EN & SRAM_DATA_EN;
    --Constants
    SRAM_CE_N <= '0';
    SRAM_UB_N <= '0';
	SRAM_LB_N <= '0';
	--Always driving SRAM_DQ unless WE
	SRAM_OE_N <= '0';
	--SRAM_DQ to IO_BUS
	IO_BUS: LPM_BUSTRI
	GENERIC MAP (
		lpm_width => 16
	)
	PORT MAP (
		data     => SRAM_DQ,
		enabledt => SRAM_DATA_EN AND IO_CYCLE,
		tridata  => IO_DATA
	);
	--SRAM_DATA to SRAM_DQ
	IO_SRAM: LPM_BUSTRI
	GENERIC MAP (
		lpm_width => 16
	)
	PORT MAP (
		data     => SRAM_DATA,
		enabledt => IO_DATA_INT,
		tridata  => SRAM_DQ
	);

	--State machine
    PROCESS(CLOCK, RESETN)
      BEGIN
        IF RESETN = '0' THEN
          STATE <= IDLE;
        ELSIF (RISING_EDGE(CLOCK)) THEN
		  CASE STATE IS
            WHEN IDLE =>
              SRAM_WE_N <= '1';
              IO_DATA_INT <= '0';
			  CASE SRAM_MODE IS
				WHEN "1100" => STATE <= SET_HIGH;
				WHEN "1010" => STATE <= SET_LOW;
				WHEN "1001" => STATE <= WRITE_DATA;
				WHEN OTHERS => STATE <= IDLE;
			  END CASE;
			WHEN SET_HIGH =>
			  SRAM_ADDR(17 DOWNTO 16) <= IO_DATA(1 DOWNTO 0);
			  CASE SRAM_MODE IS
				WHEN "1100" => STATE <= SET_HIGH;
				WHEN OTHERS => STATE <= IDLE;
			  END CASE;
			WHEN SET_LOW =>
			  SRAM_ADDR(15 DOWNTO 0) <= IO_DATA(15 DOWNTO 0);
			  CASE SRAM_MODE IS
				WHEN "1010" => STATE <= SET_LOW;
				WHEN OTHERS => STATE <= IDLE;
			  END CASE;
			WHEN WRITE_DATA =>
			  SRAM_DATA <= IO_DATA;
			  SRAM_WE_N <= '1';
			  IO_DATA_INT <= '1';
			  STATE <= WRITE_DATA2;
			WHEN WRITE_DATA2 =>
				SRAM_WE_N <= '0';
				STATE <= IDLE;
			WHEN OTHERS =>
			  STATE <=IDLE;
          END CASE;
        END IF;
      END PROCESS;
  END a;
